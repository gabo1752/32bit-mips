module test ();
    initial
        begin
            $display("Hello!");
            $finish;
        end
endmodule